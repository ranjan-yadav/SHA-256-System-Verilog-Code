module test;
reg clk,reset;
reg [255:0]input_data;

wire [255:0]out_data;

sha_256 block(input_data,out_data,clk,reset);
initial
clk = 1'b0;
always
#750 clk = ~clk;

initial
begin
reset = 1'b0;
input_data = 255'b01100001_01100010_01100011_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010;

#1500
reset <= 1'b1;
input_data = 255'b01100001_01100010_01100011_01100100_01100101_01100110_01100111_01101000_01101001_01101010_01101011_01101100_01101101_01101110_01101111_01110000_01110001_01110010_01110011_01110100_01110101_01110110_01110111_01111000_01111001_01111010_01100001_01100010_01100011_01100100_01100101_01100110;

#1500
input_data = 255'b01100001_01100010_01100011_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010_01100010;

end

initial
#6750 $finish;

endmodule
